/***************************************************************************************************
 * Module: LCMS2012_xem6010_top
 *
 * Description: This top module is for use with the Opal Kelly XEM6010 board.
 *
 * Created: Fri 22 Jul 2011 14:05:17 EDT
 *
 * Author:  Berin Martini // berin.martini@gmail.com
 **************************************************************************************************/
`ifndef _xem6010_template_ `define _xem6010_template_


`timescale 1ns / 1ps

//`include "LCMS2010_project.v"
//`include "okLibrary.v"


module LCMS2012_xem6010_top(
	input  [7:0]		hi_in,
	output [1:0]		hi_out,
	inout  [15:0]		hi_inout,
	inout					hi_aa,
	output				hi_muxsel,
//	input					reset,

	output				i2c_scl,
	output				i2c_sda,

	input					PLL_CLK1,					//PLL_CLK1 is from the PLL, expected to be 100 MHz
	input					PLL_CLK2,					//PLL_CLK2 is from the PLL, expected to be 20 MHz (for the ADC)
	output  [7:0]		LED,
	output				INT_CAPSELECT1,
	output				INT_CAPSELECT2,
	output				RES_SELECT,
	output				POST_CAPSELECT,
	output				POST_BYPASS,
	output				LPF_BYPASS,	 
	output				CDS_BYPASS,
	output				CDS_CLK1,
	output				CDS_CLK2,
	output				INFILTER_SELN,
	output				ADDR0,
	output				ADDR1,
	output				ADDR2,	 
	output				ADDR3,	 
	output 				INT_RESET,		
	output 				POST_RESET,
	output				DAC_SCLK,
	output				DAC1_SYNC,
	output				DAC2_DIN,
	output				DAC1_DIN,
	output				DAC2_SYNC,
	output				ADC_SDI,	
	output				ADC_SCK,
	output				ADC_CNV,
	input					ADC_SDO,
	output				ADC_CNV_START,  //for debug, delayed version of ADC_FS_PULSE
	output				DAC_START,		 //for debug
	output				ADC_FS_PULSE	 //for debug
	//	output [0:28] xbusp,
	//	output [0:28] xbusn,
	//	output [0:28] ybusp,	
	//	output [0:28] ybusn
	);


	/************************************************************************************
	* Internal signals
	************************************************************************************/
	localparam NUM_WIRE_IN      = 21; // start addr 8'h00, range 0 - 31,  //1 is used for the piping stuff, 19 are used for LCMS_Configuration
	localparam NUM_WIRE_OUT     = 5; // start addr 8'h20, range 0 - 31  //2 for piping stuff, 1 for adc_result_out
	localparam NUM_TRIG_IN      = 0; // start addr 8'h40, range 0 - 31
	localparam NUM_TRIG_OUT     = 0; // start addr 8'h60, range 0 - 31
	localparam NUM_PIPE_IN      = 2; // start addr 8'h80, range 0 - 31
	localparam NUM_PIPE_OUT     = 2; // start addr 8'hA0, range 0 - 31
	localparam NUM_OR           = (NUM_WIRE_OUT + NUM_TRIG_OUT + NUM_PIPE_IN + NUM_PIPE_OUT);


	// Host interface connections
	wire                    ti_clk;
	wire [30:0]             ok1;
	wire [16:0]             ok2;

	wire [(17*NUM_OR)-1:0]  ok2x;

	wire [15:0]             epWireIn    [0:31];
	wire [15:0]             epWireOut   [0:31];

	wire [0:31]             trigInClk;
	wire [0:31]             trigOutClk;
	wire [15:0]             epTrigIn    [0:31];
	wire [15:0]             epTrigOut   [0:31];

	wire [0:31]             epPipeInEn;
	wire [0:31]             epPipeOutEn;
	wire [15:0]             epPipeInData    [0:31];
	wire [15:0]             epPipeOutData   [0:31];

	//wire [7:0]              a_led;

	wire                    dcm_locked_out;
	wire                    sdram_clk;
	// synthesis attribute KEEP of sdram_clk is "true";

	wire reset;

	//clocks generated by clock divider from PLL Clock
	reg clk_1H;							//clk will be generated as 1 Hz (1 s) from the 100 MHz PLL Clock (PLL_CLK1)
	reg [27:0] clk_1H_counter;		//clk counter will be 20'h7A11F, to toggle clk every 1 s
	reg clk_1M;							//clk will be generated as 1 MHz (1 us) from the 100 MHz PLL Clock (PLL_CLK1)
	reg [15:0] clk_1M_counter;		//clk counter will be 49, to toggle clk every 1 us
	reg clk_10M;						//100 ns for now, 10 MHz
	reg [15:0] clk_10M_counter;	//dac clk counter will be 9, to toggle clk ever 10us
	

	wire [15:0] adc_result;

	LCMS2012_project #(
		.MEM_ADDR_WIDTH (10)) // # of buffer addr bits
	project (
		.a_led						(LED),

		.s_clk						(PLL_CLK1), //from PLL, 100Mhz
	//	.a_rst_hard					(reset),

		.ti_clk						(ti_clk), //opal kelly clock
		.ti_rst_soft				(epWireIn[0][0]),

		.ti_in_available			(epWireOut[0]),
		.ti_in_data_en				(epPipeInEn[0]),
		.ti_in_data					(epPipeInData[0]),

		.ti_out_available			(epWireOut[1]),
		.ti_out_data_en			(epPipeOutEn[0]),
		.ti_out_data				(epPipeOutData[0]),

		//.ti_in_test_en				(epPipeInEn[1]),
		//.ti_in_test					(epPipeInData[1]),
		//.ti_out_test_en			(epPipeOutEn[1]),
		//.ti_out_test				(epPipeOutData[1]),
		
		//signals for LCMS_configuration, signals in all caps go to the PCB (ucf connections)
		.config_clk					(clk_1M),	//1 MHz clock, to be used by LCMS configuration
		.dac_sm_clk					(clk_10M),	//clock for DAC state machine, 10 MHz
		.adc_sm_clk					(PLL_CLK2), //clock for ADC, 20 MHz
		.reset_gen_clk				(clk_1M),	//clock for the reset geberator, 1 MHz since everything here is set in us
		.reset						(reset),	
		.DAC_SCLK					(DAC_SCLK),
		.DAC1_SYNC					(DAC1_SYNC),
		.DAC1_DIN					(DAC1_DIN),
		.DAC2_SYNC					(DAC2_SYNC),
		.DAC2_DIN					(DAC2_DIN),
		.ADC_SDI						(ADC_SDI),
		.ADC_SCK						(ADC_SCK),
		.ADC_CNV						(ADC_CNV),
		.ADC_SDO						(ADC_SDO),
		.ADDR0						(ADDR0),
		.ADDR1						(ADDR1),
		.ADDR2						(ADDR2),
		.ADDR3						(ADDR3),
		.INT_CAPSELECT1			(INT_CAPSELECT1),
		.INT_CAPSELECT2			(INT_CAPSELECT2),
		.RES_SELECT					(RES_SELECT),
		.INT_RESET					(INT_RESET),
		.POST_CAPSELECT			(POST_CAPSELECT),
		.POST_RESET					(POST_RESET),
		.POST_BYPASS				(POST_BYPASS),
		.LPF_BYPASS					(LPF_BYPASS),
		.CDS_BYPASS					(CDS_BYPASS),
		.CDS_CLK1					(CDS_CLK1),
		.CDS_CLK2					(CDS_CLK2),
		.INFILTER_SELN				(INFILTER_SELN),
		//.reset						(epWireIn[1][0]),
		.addr0_i						(epWireIn[1][1]),
		.addr1_i						(epWireIn[1][2]),
		.addr2_i						(epWireIn[1][3]),
		.addr3_i						(epWireIn[1][4]),
		.int_capselect1_i			(epWireIn[1][5]),
		.post_capselect_i			(epWireIn[1][6]),
		.post_bypass_i				(epWireIn[1][7]),
		.lpf_bypass_i				(epWireIn[1][8]),
		.mode_i						(epWireIn[1][9]),		
		.int_capselect2_i			(epWireIn[1][10]),
		.res_select_i				(epWireIn[1][11]),
		.cds_bypass_i				(epWireIn[1][12]),
		.infilter_seln_i			(epWireIn[1][13]),
		.mode2_i						(epWireIn[1][14]),
		.int_gbt_i					(epWireIn[2]),
		.int_vbn_i					(epWireIn[3]),
		.int_vbp_i					(epWireIn[4]),
		.post_gbt_i					(epWireIn[5]),
		.post_vbn_i					(epWireIn[6]),
		.post_vbp_i					(epWireIn[7]),
		.obuff_gbt_i				(epWireIn[8]),
		.obuff_vbn_i				(epWireIn[9]),
		.obuff_vbp_i				(epWireIn[10]), //0A
		.vref_i						(epWireIn[11]), //0B
		//.VCMD							(epWireIn[12]), //0C   //now VCMD comes from a pipe in, not from a wire
		.reset_period_i			(epWireIn[13]), //0D
		.int_reset_duration_i	(epWireIn[14]), //0E
		.post_reset_duration_i	(epWireIn[15]), //0F
		.v_sampling_period_i		(epWireIn[16]), //10    //wireIn is available from 00 up to 1F (32 wireIns total)
		.adc_result					(adc_result[15:0]),
		.start_meas					(epWireIn[17][0]), //11  start is bit 0 of wirein 17, or it could be moved to wire in 1 bit 10
		.cds_time1_delay_i		(epWireIn[18]), //12
		.cds_time2_delay_i		(epWireIn[19]), //13
		.cds_width_i				(epWireIn[20]), //14
		.adc_cnv_start				(ADC_CNV_START),  //only output this for debug, generated within lcms2012_project
		.dac_start					(DAC_START),      //only output this for debug, generated within lcms2012_project
		.adc_fs_pulse				(ADC_FS_PULSE)		//only output this for debug, generated within lcms2012_project, delayed version of ADC_CNV_START
		);


    /************************************************************************************
     * Instantiate the Opal Kelly okHost and okWireOR, connect endpoints
     ************************************************************************************/

    assign hi_muxsel = 1'b0;

    okHost
    okHI (
        .hi_in      (hi_in),
        .hi_out     (hi_out),
        .hi_inout   (hi_inout),
        .hi_aa      (hi_aa),
        .ti_clk     (ti_clk),
        .ok1        (ok1),
        .ok2        (ok2) );


    okWireOR #(.N(NUM_OR)) wireOR (ok2, ok2x);


    genvar wi;
    generate
        for (wi = 0; wi < NUM_WIRE_IN; wi = wi + 1) begin: WI_

            okWireIn
            wire_in (
                .ok1        (ok1),
                .ep_addr    (8'h00 + wi),
                .ep_dataout (epWireIn[wi]) );

        end
    endgenerate


    genvar wo;
    generate
        for (wo = 0; wo < NUM_WIRE_OUT; wo = wo + 1) begin: WO_

            okWireOut
            wire_out (
                .ok1        (ok1),
                .ok2        (ok2x[wo*17 +: 17]),
                .ep_addr    (8'h20 + wo),
                .ep_datain  (epWireOut[wo]) );

        end
    endgenerate


    genvar ti;
    generate
        for (ti = 0; ti < NUM_TRIG_IN; ti = ti + 1) begin: TI_

            okTriggerIn
            trigger_in (
                .ok1        (ok1),
                .ep_addr    (8'h40 + ti),
                .ep_clk     (trigInClk[ti]),
                .ep_trigger (epTrigIn[ti]) );

        end
    endgenerate


    genvar to;
    generate
        for (to = 0; to < NUM_TRIG_OUT; to = to + 1) begin: TO_

            okTriggerOut
            trigger_out (
                .ok1        (ok1),
                .ok2        (ok2x[(NUM_WIRE_OUT+to)*17 +: 17]),
                .ep_addr    (8'h60 + to),
                .ep_clk     (trigOutClk[to]),
                .ep_trigger (epTrigOut[to]) );

        end
    endgenerate


    genvar pi;
    generate
        for (pi = 0; pi < NUM_PIPE_IN; pi = pi + 1) begin: PI_

            okPipeIn
            pipe_in (
                .ok1        (ok1),
                .ok2        (ok2x[(NUM_WIRE_OUT+NUM_TRIG_OUT+pi)*17 +: 17]),
                .ep_addr    (8'h80 + pi),
                .ep_write   (epPipeInEn[pi]),
                .ep_dataout (epPipeInData[pi]) );

        end
    endgenerate


    genvar po;
    generate
        for (po = 0; po < NUM_PIPE_OUT; po = po + 1) begin: PO_

            okPipeOut
            pipe_out (
                .ok1        (ok1),
                .ok2        (ok2x[(NUM_WIRE_OUT+NUM_TRIG_OUT+NUM_PIPE_IN+po)*17 +: 17]),
                .ep_addr    (8'hA0 + po),
                .ep_read    (epPipeOutEn[po]),
                .ep_datain  (epPipeOutData[po]));

        end
    endgenerate

	/************************************************************************************
	* Implementation
	************************************************************************************/

	assign i2c_scl  = 1'bz;
	assign i2c_sda  = 1'bz;
	
	assign reset = epWireIn[1][0];	
	//reg [7:0] msb;
	//assign led = adc_result[15:8];
	//	reg [7:0] lsb;
	assign epWireOut[2] = {adc_result[15:0]};
	assign epWireOut[3] = {epWireIn[16][15:0]};
	//assign epWireOut[2][15:0] = {adc_result[15:0]};
	//assign epWireOut[3] = {adc_result[15:0]};
	//assign epWireOut[2] = {adc_result[15:8], 8'b11111111};
	//assign epWireOut[3] = {adc_result[7:0]};
	
//	reg a;
	
//	always @ (posedge clk_1H, posedge reset) begin
//		if (reset) begin
//			a <= 0;
//		end
//		else begin
//			a <= !a;
//			if (a) msb = adc_result[15:8];
//			else	 msb = adc_result[7:0];
//		end
//	end
	
	//generate a slow 1s clock signal so we can control stuff
//	always @ (posedge PLL_CLK1, posedge reset) begin
//		if (reset) begin
//			clk_1H_counter <= 0;
//			clk_1H <= 0;
//		end
//		else begin	
//			clk_1H_counter <= clk_1H_counter + 1'b1;
//			if (clk_1H_counter == 28'h2FAF07F) begin
//				clk_1H_counter <= 28'h0000000;
//				clk_1H <= !clk_1H;
//			end
//		end
//	end	
	
	//generate 1 MHz (1 us) clock signal from input 100MHz PLL_CLK1 pll
	always @ (posedge PLL_CLK1, posedge reset) begin
		if (reset) begin
			clk_1M_counter <= 0;
			clk_1M <= 0;
		end
		else begin	
			clk_1M_counter <= clk_1M_counter + 1'b1;
			if (clk_1M_counter == 16'D49) begin
				clk_1M_counter <= 16'D0;
				clk_1M <= !clk_1M;
			end
		end
	end
	
	
	//generate 10 MHz (100 ns) clock signal from input 100MHz PLL_CLK1 pll
	always @ (posedge PLL_CLK1, posedge reset) begin
		if (reset) begin
			clk_10M_counter <= 0;
			clk_10M <= 0;
		end
		else begin	
			clk_10M_counter <= clk_10M_counter + 1'b1;
			if (clk_10M_counter == 16'D4) begin
				clk_10M_counter <= 16'D0;
				clk_10M <= !clk_10M;
			end
		end
	end
	
	// old stuff from Berin
	    assign trigInClk[0]     = ti_clk;
	    assign trigOutClk[0]    = ti_clk;

	//    assign led      = ~{a_led, dcm_locked_out};
		
		
//		assign led = 8'b0;
//		assign INT_CAPSELECT = 1'b1;
//		assign POST_CAPSELECT = 1'b1;
//		assign POST_BYPASS = 1'b1;
//		assign LPF_BYPASS = 1'b1;
//		assign ADDR0 = 1'b1;
//		assign ADDR1 = 1'b1;
//		assign ADDR2 = 1'b1;
//		assign ADDR3 = 1'b1;
//		assign DAC_SCLK = 1'b1;
//		assign DAC1_SYNC = 1'b1;
//		assign DAC2_DIN = 1'b1;
//		assign DAC1_DIN = 1'b1;
//		assign DAC2_SYNC = 1'b1;
//		assign ADC_SDI = 1'b1;
//		assign ADC_SCK = 1'b1;
//		assign ADC_CNV = 1'b1;
//		assign ADC_SDO = 1'b1;
		
//		assign led[0] = reset;
//		assign led[1] = PLL_CLK1;
//		assign led[2] = clk;
//		assign led[3] = 1'b1;
//		assign led[4] = 1'b1;
//		assign led[5] = 1'b1;
//		assign led[6] = 1'b1;
//		assign led[7] = 1'b1;
//		
//		assign xbusp[0]= 1'b1;
//		assign xbusp[1]= 1'b1;
//		assign xbusp[2]= 1'b1;
//		assign xbusp[3]= 1'b1;
//		assign xbusp[4]= 1'b1;
//
//		assign xbusp[7]= 1'b1;
//		assign xbusp[8]= 1'b1;
//		assign xbusp[9]= 1'b1;
//		assign xbusp[10]= 1'b1;
//		assign xbusp[11]= 1'b1;
//		assign xbusp[12]= 1'b1;
//		assign xbusp[13]= 1'b1;
//		assign xbusp[14]= 1'b1;
//		assign xbusp[15]= 1'b1;
//		assign xbusp[16]= 1'b1;
//		assign xbusp[17]= 1'b1;
//		assign xbusp[18]= 1'b1;
//		assign xbusp[19]= 1'b1;
//		assign xbusp[20]= 1'b1;
//		assign xbusp[21]= 1'b1;
//		assign xbusp[22]= 1'b1;
//		assign xbusp[23]= 1'b1;
//		assign xbusp[24]= 1'b1;
//		assign xbusp[25]= 1'b1;
//		assign xbusp[26]= 1'b1;
//		assign xbusp[27]= 1'b1;
//		assign xbusp[28]= 1'b1;
//
//		assign xbusn[0]= 1'b1;
//		assign xbusn[1]= 1'b1;
//		assign xbusn[2]= 1'b1;
//		assign xbusn[3]= 1'b1;
//		assign xbusn[4]= 1'b1;
//		assign xbusn[5]= 1'b1;
//		assign xbusn[6]= 1'b1;
//		assign xbusn[7]= 1'b1;
//		assign xbusn[8]= 1'b1;		
//		assign xbusn[9]= 1'b1;
//		assign xbusn[10]= 1'b1;
//		assign xbusn[11]= 1'b1;
//		assign xbusn[12]= 1'b1;
//		assign xbusn[13]= 1'b1;
//		assign xbusn[14]= 1'b1;
//		assign xbusn[15]= 1'b1;
//		assign xbusn[16]= 1'b1;
//		assign xbusn[17]= 1'b1;
//		assign xbusn[18]= 1'b1;
//		assign xbusn[19]= 1'b1;
//		assign xbusn[20]= 1'b1;
//		assign xbusn[21]= 1'b1;
//		assign xbusn[22]= 1'b1;
//		assign xbusn[23]= 1'b1;
//		assign xbusn[24]= 1'b1;
//		assign xbusn[25]= 1'b1;
//		assign xbusn[26]= 1'b1;
//		assign xbusn[27]= 1'b1;
//		assign xbusn[28]= 1'b1;
//		
//		assign ybusp[0]= 1'b1;
//		assign ybusp[1]= 1'b1;
//		assign ybusp[2]= 1'b1;
//		assign ybusp[3]= 1'b1;
//		assign ybusp[4]= 1'b1;
//		
//		assign ybusp[7]= 1'b1;
//		assign ybusp[8]= 1'b1;
//		assign ybusp[9]= 1'b1;
//		assign ybusp[10]= 1'b1;
//		assign ybusp[11]= 1'b1;
//		assign ybusp[12]= 1'b1;
//		assign ybusp[13]= 1'b1;
//		assign ybusp[14]= 1'b1;
//		assign ybusp[15]= 1'b1;
//		assign ybusp[16]= 1'b1;
//		assign ybusp[17]= 1'b1;
//		assign ybusp[18]= 1'b1;
//		assign ybusp[19]= 1'b1;
//		assign ybusp[20]= 1'b1;
//		assign ybusp[21]= 1'b1;
//		assign ybusp[22]= 1'b1;
//		assign ybusp[23]= 1'b1;
//		assign ybusp[24]= 1'b1;
//		assign ybusp[25]= 1'b1;
//		assign ybusp[26]= 1'b1;
//		assign ybusp[27]= 1'b1;
//		assign ybusp[28]= 1'b1;
//		
//		assign ybusn[0]= 1'b1;
//		assign ybusn[1]= 1'b1;
//		assign ybusn[2]= 1'b1;
//		assign ybusn[3]= 1'b1;
//		assign ybusn[4]= 1'b1;
//		assign ybusn[5]= 1'b1;
//		assign ybusn[6]= 1'b1;
//		assign ybusn[7]= 1'b1;
//		assign ybusn[8]= 1'b1;
//		assign ybusn[9]= 1'b1;
//		assign ybusn[10]= 1'b1;
//		assign ybusn[11]= 1'b1;
//		assign ybusn[12]= 1'b1;
//		assign ybusn[13]= 1'b1;
//		assign ybusn[14]= 1'b1;
//		assign ybusn[15]= 1'b1;
//		assign ybusn[16]= 1'b1;
//		assign ybusn[17]= 1'b1;
//		assign ybusn[18]= 1'b1;
//		assign ybusn[19]= 1'b1;
//		assign ybusn[20]= 1'b1;
//		assign ybusn[21]= 1'b1;
//		assign ybusn[22]= 1'b1;
//		assign ybusn[23]= 1'b1;
//		assign ybusn[24]= 1'b1;
//		assign ybusn[25]= 1'b1;
//		assign ybusn[26]= 1'b1;
//		assign ybusn[27]= 1'b1;
//		assign ybusn[28]= 1'b1;


endmodule

`endif //  `ifndef _xem6010_template_
